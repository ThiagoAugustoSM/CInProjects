module projetoGeral(
	IorD,
	WR,
	AluSrcA,
	AluSrcB,
	AluOP,
	PCsrc,
	PCwrite,
	IRwrite,
	muxR1
);



endmodule
