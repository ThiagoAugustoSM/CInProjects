module mux();